library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Funkcja_f_tablica_vhdl is
    Port ( w, x, y, z : in  STD_LOGIC;
           f : out  STD_LOGIC);
end Funkcja_f_tablica_vhdl;

architecture Behavioral of Funkcja_f_tablica_vhdl is

begin



end Behavioral;

